module QR;initial begin $write("%s",("let s=(\"Module QR\\n\")\nput=s\nprint\nlet s=(\"Sub Main()\\n\")\nput=s\nprint\nlet s=(\"Dim c,n:Dim s As Object=System.Console.OpenStandardOutput():Dim t()As Short={26,34,86,127,148,158,200}:For Each d in\\\"BasmCBBBCRE`F<<<<C<`C<B`BBD#CXwasi_snapshot_preview1Jfd_writeBBEEDCDGECB@IUDHmemoryDBH_startBDL|DRBAC BAJlACA4RB9MiCD<AERCA>D!BE@ABRCABRCABRCAJ!CE@ B-BB CACk:CvACqRC COBMADRCACRCADRCABRCABRC BACj:B-BBOBMADRCADRCADRCAFRCMM}CBABM~(BBBCBBB,BBBDBBB0BBBDBBB4BBB=BBB?BBB;BBB ...\\\\t..\\\\n..(module(import :wasi_snapshot_preview1: :fd_write: (func(param i32 i32 i32 i32)(result i32)))(memory(export :memory:)(data :\\\\08\\\\00\\\\00\\\\00$:))(func(export :_start:)i32.const 1 i32.const 0 i32.const 1 i32.const 0 call 0 drop))\\\":c=Asc(d):If c=36:For c=0To 11:s.WriteByte(If(c Mod 3,Asc(6"));
$write("%s",("23475.ToString(\\\"x8\\\")(1Xor 7-c*2\\\\3)),92)):Next:Else:n=(c>124)*(8*c-40261):Do While n>127:s.WriteByte(128+(127And n)):n\\\\=128:Loop:s.WriteByte(If(c<125,If((c-1)\\\\7-8,c+66*(c>65And c<91),t(c-57)),n)):End If:Next:For Each c in\\\"<?xml version='1.0'?><?xml-stylesheet type='text/xsl'href='QR.xslt'?><xsl:stylesheet version='1.0' xmlns:xsl='http://www.w3.org/1999/XSL/Transform'><xsl:output method='text'/><xsl:template match='/'><![CDATA[sub f(s$,n)print(s$);:for i=1to n print(\\\"\\\"\\\\\\\\\\\"\\\");:next:end sub:f(\\\"\\\"write,format=\\\\\\\"\\\"%s%s%s%s\\\\\\\"\\\",\\\\n(\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"write{-}{txt}{echo -E $'(\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\"with Ada.Text_Io;procedure qr is begin Ada.Text_Io.Put(\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans B(Buffer)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f("));
$write("%s",("\\\"\\\"\\\\\\\"\\\"trans O(n)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"B:add(Byte(+ 128 n))\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans f(v n)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(+(/ n 64)107)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(n:mod 64)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O v\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans D(n)\\\"\\\",2):f(\\\"\\\"{if(< n 4)\\\"\\\",2):f(\\\"\\\"{f(+(* 6 n)9)48\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{if(n:odd-p)\\\"\\\",2):f(\\\"\\\"{D(- n 3)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9"));
$write("%s",("):f(\\\"\\\"\\\\\\\"\\\"f 27 48\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 36 11\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{D(/ n 2)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 21 48\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 48 20\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans S(Buffer\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"STRINGz:=REPR226+REPR153,a:=z+REPR166,b:=a+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"2\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR160,c:=b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR165,t:=\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class QR\\\"\\\",2"));
$write("%s",("):f(\\\"\\\"{public static void main(String[]a)\\\"\\\",2):f(\\\"\\\"{a=(\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"write(\\\"\\\",4):f(\\\"\\\"'implement main0()=print(^1^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"BEGIN\\\"\\\",2):f(\\\"\\\"{print(^3^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"echo ^1^\\\"\\\",4):f(\\\"\\\"'f(s)\\\"\\\",2):f(\\\"\\\"{System.out.print(s);\\\"\\\",2):f(\\\"\\\"}s=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"389**6+44*6+00p45*,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(c:(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"#include<stdio.h>^8^"));
$write("%s",("nchar*p=(^15^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Ra#include<iostream>^16^nint main()\\\"\\\",2):f(\\\"\\\"{std::cout<<(^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class Program\\\"\\\",2):f(\\\"\\\"{public static void M83abbSystem.Console.Write(^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Quine Relay Coffee.^64^n^64^nIngredients.^64^n^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");for(int i=9;i++<126;)[3pva$^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"} g caffeine \\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"}I3b54rja^64^nMethodv4f#aeach(char c in(^6"));
$write("%s",("3^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")))^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2al3dp3c[2cs3c,3l[2k@3kqa^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")s rts(ecalper.h3eja^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"     53c4a SUTATS(egassem^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"rts(nltnirp(])]^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NUR POTSu4cba.C3dh3dX3bba[65bX4df5lp3lna\\\"\\\",2):f(\\\"\\\"})1(f\\\"\\\",2"));
$write("%s",("):f(\\\"\\\"{#\\\"\\\",2):f(\\\"\\\"};)06xt3ciaqp]^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'[p]13nfa3(f\\\"\\\",2):f(\\\"\\\"{#w3nga7(f\\\"\\\",2):f(\\\"\\\"{#.x3nga51(f\\\"\\\",2):f(\\\"\\\"{##4nM3sca3643qw3yf6dx3kca\\\"\\\",2):f(\\\"\\\"};l4tda,43z3sma^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\""));
$write("%s",(",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' D ; EYB RCc4tC3pka721(f\\\"\\\",2):f(\\\"\\\"{#DNE;34da. A\\\"\\\",2):f(\\\"\\\"{47eaPOTS|48\\\"\\\",2):f(\\\"\\\"{45oaRQ margorp dneF34baS^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'46%8-ca83737ba&J4-93bgaS POOLv87ba^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'83[83ida&,)-96ga. TNUO655fa(rahcX6.%4dgaB OD 0096ca&,\\\"\\\",2):f(\\\"\\\"{83ca)AW87R86qaEUNITNOC  "));
$write("%s",("    01)66~67D5/n>deaRC .>34ka,1=I 01 OD[@8caPU?35)83va;TIUQ;)s(maertSesolC;XHeN3$ra598(f\\\"\\\",2):f(\\\"\\\"{#tiuqn\\\"\\\",2):f(\\\"\\\"})420:41pa9191(f\\\"\\\",2):f(\\\"\\\"{#n\\\"\\\",2):f(\\\"\\\"})84022HxX5qca69mIy[Grca08<H3ea5526~A[83odamifR4.fa93623R4[83nbatN45%a315133A71/129@31916G21661421553/Y35wa%%%%\\\"\\\",2):f(\\\"\\\"}*+1%%%%811 -\\\"\\\",2):f(\\\"\\\"})867\\\"\\\",2):f(\\\"\\\"{3ahaj:+1 j@a45baw:35935baW:35ba\\\"\\\",2):f(\\\"\\\"{:35va)(esolc.z;)][etyb sa):9[83;ea9746(?au4[83jba,t4[83jea!\\\"\\\",2):f(\\\"\\\"})8j3aca~~#4[83jea(rt.w4[83jba)<5eda\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};m3ffa~~dnep3ira~~~~PUEVIGESAELPnr3ala~~1,TUODAERw3a73k$a(etirw;\\\"\\\",2):f(\\\"\\\"};u=:c;))652%%%%)u-c((||23kda#-<r3kda||i+3nhaBUS1,ODw4rka)3/4%%%%i(S4c~5l[4yPa2=:/t;2%%%%t+2*u=:u\\\"\\\",2):f(\\\"\\\"{od7 ot0 yreve;i-=:u;1=:+i\\\"\\\",2):f(\\\"\\\"{od))1(ev"));
$write("%s",("om(dro=:t elihw?s;)s*:5pm5ww3kn7dladohtem dne.s3dganrutern3d~aV);gnirtS/gnal/avajL(nltnirp/GKa|atnirP/oi/avaj lautrivekovniJ3d/4k[2cib\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};0=q;)]q[c=z(tnirp.tuo.metsyS;)0(tArahc.y+z=]++n[c;y:]q[c?n<q=y\\\"\\\",2):f(\\\"\\\"{)0>2%%%%++i(fi;48%%%%)31-)i>3c&as(+87*q=q\\\"\\\",2):f(\\\"\\\"{);41712<i;(rof;n)rahc(+L4s[2k+3^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'oa=]n[c);621<n++t4aqa0=q,0=n,0=i tni;O3^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\""));
$write("%s",("\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'Ub6a5k4asdRbQexmxf\\\"\\\",2):f(\\\"\\\"}hpm0g<bedRb;fW-;agb-a|dzdxd0gGb8aqeRdYd5a,LUi;agb-epb>aqeRddgJaBd8gFbaeIfOa5aacLipY6f9aKu4aLa7a;a\\\"\\\",2):f(\\\"\\\"}|5a33kdxd;aNa?c6a|eebHaFaIaebzeJaeb9a/a6a2dQbUe-f2a-E3cdacEeC3g/a-f/aof0f0gH55aDm.b2e6aRa;dJZzgPa1bli;aTapc?3a6b5kof6amc<b-a6a-fYmsbYg.2Ii4atcSiU2tkWYtkYR\\\"\\\",2):f(\\\"\\\"}bJaMa\\\"\\\",2):f(\\\"\\\"}bUbtk9sJaJaUa-bJaMdJa8bKX;a8bG-Ka8bG-8be@kCPaOaX9NaT=Ka;1BJTa8b*\\\"\\\",2):f(\\\"\\\"{G-8bU2wb\\\"\\\",2):f(\\\"\\\"}bJaLaJa8b*\\\"\\\",2):f(\\\"\\\"{U2j4c\\\"\\\",2):f(\\\"\\\"{a8bU24bU2:b+bWYtkWYwbkCJaHa\\\"\\\",2):f(\\\"\\\"{3a;3ajbHaJaFdc\\\"\\\",2):f(\\\"\\\"{;a;1Ua:aUa:aKXyhycwh>athAa2aUe?a7a6a=g:a?aMboh6a?e:a*02a?a1a,hMbogiihhKg,nIfbh4aqqsbsb2be3^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\""));
$write("%s",("\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'+ayhDa-a.2WgQbwg<b=a-a6l*c3bxdUe=aJg+<9ag3cra2bMa7a=h;h9h7h5h9k3f?aAdb6Pcgfvftioi7a<h?l=lMa6l*cEc,dJa>a2aIf;f9fMa?a+<Hi/i-i6a/3iUaxdtbA*-i/aTh=a;i.\\\"\\\",2):f(\\\"\\\"}-c.\\\"\\\",2):f(\\\"\\\"}OaqFi,Na;i=k6a7bem0gwblkUe2b5ax2Gj4b-bhc,oxkxk|oPfxd;aaiXj3;aea6a2bc;egc1CvY6aAo2a5a3a@Q\\\"\\\",2):f(\\\"\\\"{kobRl6uxk6azi|oHa:eelcm;a|mQaw/0gLM<b3bxd6aniKl5a6jAV6i\\\"\\\",2):f(\\\"\\\"}h\\\"\\\",2):f(\\\"\\\"{hPa;aFjcc8bfbpbK;*wZbfynb\\\"\\\",2):f(\\\"\\\"{gdkbk4i,7FldlwlFm<b<b<bIk:b@k<b<b,cNkKk7b-bNkEaKo3bDd7lul9atqSf5bC\\\"\\\",2):f(\\\"\\\"},cNk=a9a7bubq3emaEaNl9l,cNkAa/3aeaeM8f=3a-3ieaJbupM3g#aDaCaBa>a9a7bwbSfeMr4+lYjJl,cNki3a)a+n3"));
$write("%s",("h.b1h,cNksb0g?a@jkmagimZkGkEa3a6as3eqajl6aelcmul5l<bzeG?e^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3eeaAl3a)3coaFOBG\\\"\\\",2):f(\\\"\\\"}W0cDm*kBm^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3ewaOlrh6a<b6iLj?Q2b2a2aH6/3aWabMLf4gwblk0g@a>anc:e7b5aIi=anbggyb/l5a,bJa6a-bJaJaubXh;dHawblkHa:e-b9a9b9aAl5aigshm3atb@a8eig6a@a>a:a|b9a0b9a@a>a7a6a@a>e|b5a:a9bJa0b5aig6a-b9aAl9aN=Ja9bggnbJa6a|b5a,b0g:e-b5a>O-a5h9apb6ky"));
$write("%s",("4uYAig3draa8bAdli-aLMQ2bb-ay3eba7y3hcaLMv6ecaMl,6aj6akaXb;d9f/bxd:4a^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'a8b9a7bJcJayb>a8hGaihJa*cicfg?b,bFaq3a2a-b-a8gUe@a>aJu5aDcC::atcJaub5aEcxb,7,b4b-bJa3H8hkaamEkmdqi0gp8os3aDdgm3apb;awblk/md2BEAGFO<Sy4LKtYJdHd1m>oLM1Cy4uY:SJoRmaoDoin|nXoHoW,mI.bB79|36?6EB1YIs+\\\"\\\",2):f(\\\"\\\"{eyjbepky+l55Ssm9b-as.b\\\"\\\",2):f(\\\"\\\"{TXpCaaP/b:GypkbEalb.baDypu+qqe6-b>y1pepcWjHgb1EZahb=atc6hNGhb?aP9ibubuAYadbeb@PAaNvjbDa+Tgb61<0Na99ib=Mb-V5>qkbn\\\"\\\",2):f(\\\"\\\"},XV<Ea>r<zhbEawbuv7be<ZYQw9wRRI.lbqEOptbYZBWWa2-tbibR6j\\\"\\\",2):f(\\\"\\\"{CaaP\\\"\\\",2):f(\\\"\\\"{bYa2\\\"\\\",2):"));
$write("%s",("f(\\\"\\\"}Za.;,K|=Qxz:rsgDXxabq<\\\"\\\",2):f(\\\"\\\"{rr?B7cb8bSw6k*6a&dIDt0HuBtID,Cub@4tbYw@ayMhz+v,pf:XpKqI.Vaxbcu\\\"\\\",2):f(\\\"\\\"{ufr>anFs.L0X:L-bO*b,b;Ker+lGpDa8r.bWaubtT9bWar91u8;>a=pSad1YavbdqBsyuVaCrcbM+jBB\\\"\\\",2):f(\\\"\\\"}-b.rBp1L;:xp|,,1x\\\"\\\",2):f(\\\"\\\"{xbxbz.=aybZqjbD2<yT0upUa?1NaKqW+E\\\"\\\",2):f(\\\"\\\"}6-3=kbevPavvQPsM*bmbuphjNaDaWp4b7\\\"\\\",2):f(\\\"\\\"{uf-bmuCstD5/f?z1X*G+T48q6we@j\\\"\\\",2):f(\\\"\\\"{Wa.tm*Na8t;B3b-sibKqeMpTz\\\"\\\",2):f(\\\"\\\"{YarqA12@8+c;gMLvvCfqoxabrsC9c*dBOEy2bKqe:kb7wHJyb6bwb2bOajbDyUae;DSXa8q3ZkbK,iEQqspkr-bvp6z?\\\"\\\",2):f(\\\"\\\"}>vl1<ajb2ba?7Edbb<Ya090b6Fb<YaItj1xrOWsx=pS;.p;-7tJwD2H98+\\\"\\\",2):f(\\\"\\\"{bq.x8hbjb19D=\\\"\\\",2):f(\\\"\\\"{0jbO1AHNO<7aPeUhb6b0b9bF7.:>-m2jb.\\\"\\\",2):f(\\\"\\\"}EsJNDank.:vbPq:27E0NnWuby9=JAa-.4@jb9b,b9+l-*7\\\"\\\",2):f(\\\"\\\"{0-bar/pCrjbZap>?1lb"));
$write("%s",("DaR5:KuWl>jbDaG.DaJNDaB1*>lqe@3<SLspJN.:Qq.:wb6hf5EajbIqUngb*bY9cea6bCay3aud@T\\\"\\\",2):f(\\\"\\\"{:L-r30.;09T\\\"\\\",2):f(\\\"\\\"{:Ts,bh;/TzpLXYa0T.TSW1,*T16\\\"\\\",2):f(\\\"\\\"{TL-jbxTWayr;sh;hbiSYQzrq\\\"\\\",2):f(\\\"\\\"{spvbE.QaZqIGL-.p,CspJC.:gkTal2SajbQaLxQWVS.:GDspo7CvJSd|cpLXcbyp9ZlbAX?1;7N2.bvr+bBBK7/p/bkrTaDj|Jf5=aRwp3ubDansspkrjbDaPw.:krjbRrhzNap3ubRr*IgbS+K@/ZyS9b6<Rr\\\"\\\",2):f(\\\"\\\"}b-bJZ||DavxPaSQt0n4jsp2,bZRjq2bc>\\\"\\\",2):f(\\\"\\\"}y7bWYDawb.ZhWdpg*5A2*6dhdhqDaIpEpCa+rDaB1YqxZk,cbH2bSibOpjbyb|RuxHp4bDaNwGIHIwbhbkblRjblbhb?a3\\\"\\\",2):f(\\\"\\\"{hb?a8bhb130baEjsUX,xA=64n4-VcbmPbrhbhbDu?aZJDa13+1O+J>hbRau--0yMKZ-0yMlRzrhbRaop49XT:*1/n1\\\"\\\",2):f(\\\"\\\"{T:qk\\\"\\\",2):f(\\\"\\\"{H.DanDUxs6hbYa>a3\\\"\\\",2):f(\\\"\\\"{hbm-MGZ|N;bSYavbubQ2ub3bVvibgWzL5;.;ap4bEavpJq0pvbCvq4YaGug*f,fb>a*3efdb@a4bDL8"));
$write("%s",("bd4PaM3+>6cU3IM3aea@tAag5-fcQaZUNAiShb4\\\"\\\",2):f(\\\"\\\"}J;A?Phz\\\"\\\",2):f(\\\"\\\"{CrZtKO;pG424CrjbiDBa;Y8+*XmRhb,qAaf:\\\"\\\",2):f(\\\"\\\"{0+1\\\"\\\",2):f(\\\"\\\"{pj1*\\\"\\\",2):f(\\\"\\\"}G\\\"\\\",2):f(\\\"\\\"{>+Tz\\\"\\\",2):f(\\\"\\\"{085MpKp4b3+JZDa\\\"\\\",2):f(\\\"\\\"}+k;TaYa8bDwYaz5hzGaNZo:VB4*Xp+1\\\"\\\",2):f(\\\"\\\"{pp2hb0bYatb\\\"\\\",2):f(\\\"\\\"}b4sybLuTsW2@Asqfr+b9+vbhw=p0Y>4iHzb2@c4Aa@rvz8|:dxd2bXxydV>0lRquZvW@,sWPqV.6*g8A>*\\\"\\\",2):f(\\\"\\\"{3=nWG+vQ3b6tJQ?/LLgz>87w.>JZlbYYJS|bRC,L;0kGju4:j9ritb<5,1|rabybvbVvrsov\\\"\\\",2):f(\\\"\\\"}pFa+1rsgb*:VaEsct=Lyb|X+ba-XP:2arU5fsFag<7NCSt?mbb*LxvrMZyb\\\"\\\",2):f(\\\"\\\"}7YArqTayb0b?a;:abx2mO=Mv?Du*bej3WSa\\\"\\\",2):f(\\\"\\\"}gWuTaf-3beyhxYa130b?aQDFaXa7q14XUC7=/Mh@0p-ZaTr5bufi>c:CaMp.dKR>8ybabgM?vEqCrlEXaTO~6c-c*v*bj\\\"\\\",2):f(\\\"\\\"}Ra5,OaTa<s2KH=mx<IfHy\\\"\\\",2):f(\\\"\\\"}<6Muzg.tKsLi"));
$write("%s",(":Tbvhj2Da>C3Jsam|bj9?a|bQBCajK>K,b**.Qczt|R9-dB3vb/M7v-Mw\\\"\\\",2):f(\\\"\\\"}0qcyZ8|syjw\\\"\\\",2):f(\\\"\\\"}=a-4=R/x07zg>BTFybwb73Gv@a3bILUalv7bo|Crcbg8t+.7sICSpU/bl+UYYatb2Wts.bhbi-MSvHO02\\\"\\\",2):f(\\\"\\\"}Va?adz=Lebk-p01h-+YZz6OIa?a;sP\\\"\\\",2):f(\\\"\\\"}1rQ=*iCr8qiy1bAXU2LCIjRaLT*\\\"\\\",2):f(\\\"\\\"}XVIt9uO=iyJwF-k-tF*\\\"\\\",2):f(\\\"\\\"}x-LTRKx6c&fetnvaD1y78n*>6E|@aXa9blb3bffj.GGzb3LUTgz4EOX6p\\\"\\\",2):f(\\\"\\\"}gb95+OhN9L2dzZa/ysz\\\"\\\",2):f(\\\"\\\"{bY8:3N<k-N<hwp0*tx\\\"\\\",2):f(\\\"\\\"}/ttbmWAt*z>6\\\"\\\",2):f(\\\"\\\"}b\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"XaE0=acX*b5blHybQttbUa,\\\"\\\",2):f(\\\"\\\"}Swru9yHPj1Z;YaCa|+.7x*xbyw;3-i0vPaawaEKij.LDDaorybQaYIHt\\\"\\\",2):f(\\\"\\\"{bzvebn64bib*bp2hb8bbbzpOqC@l1PaxPVa\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{yI4b*s=a5567WBh|>-brJOb5n<Yai/5p@aNaovF@c,+bMrNq@,pTB*Eaabybh/5bnq,Vz\\\"\\\",2):f(\\\"\\\"{Lx4b*sL"));
$write("%s",("M\\\"\\\",2):f(\\\"\\\"}ABG\\\"\\\",2):f(\\\"\\\"}Wdd550wEa+luA77Vj=zvb1bVapsWBB3aJfr@x8b*b=aWakbD7d|:@Za5+dJYYrUC\\\"\\\",2):f(\\\"\\\"}Oa/uKX|9zrTv85</GaBSkb2WN|sx*bcH1b19K+PaDSw*fb3bj1hbbt*b=amU\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}UGPay9trW2x\\\"\\\",2):f(\\\"\\\"}Si-b<a53gvYaSaC/4bQtL08CCcVa#7a,bxuh|qx?a:@lb8+SiRw>=/qz|=ax577D5DSPahbFafrKu4bH1KwJx\\\"\\\",2):f(\\\"\\\"}lD7Dy<=Zl*CjbySC356VaywPWn9A*eucukyNWQavx9,W30bU3C3M\\\"\\\",2):f(\\\"\\\"{m1WaF@IG?tKO7b0Hub/1Y9ctdUaSpQRE\\\"\\\",2):f(\\\"\\\"}E\\\"\\\",2):f(\\\"\\\"{.b6bYaasL;1b*C4bGX-bVzKBQC4>ybab:\\\"\\\",2):f(\\\"\\\"{+;Ls3wQCh5tb20Wa+@b6\\\"\\\",2):f(\\\"\\\"{*VaasRRmtFrpJc:.QC5Atvuh8h5wI5blYxscpy?q.U2<7KvAa4.QzhbQ4,6<<E-MQ>Ak|f1e7evF2lEtbzgtb\\\"\\\",2):f(\\\"\\\"}bVak@vbQa,iOsiDo\\\"\\\",2):f(\\\"\\\"{QV9KlE|lX7sMOs1bjv4\\\"\\\",2):f(\\\"\\\"}i;tET\\\"\\\",2):f(\\\"\\\"{dpX\\\"\\\",2):f(\\\"\\\"}77@tJzYj8zTBlq38YakS"));
$write("%s",("IuNCDaibR72bSCN5dbCrY*TzWBB.-8>aEymHP1Epfq5bZ6J7c4*EV*q.bbq?19K9cUc/dTs>=2wo7bbUXebh8l4|bK.*=NATaZJ7bX,H,c-y/TFZUiSSG>NU02\\\"\\\",2):f(\\\"\\\"}VaAJ|7,bYAq.Sz7bSs2bmxaE1rQI;xJx\\\"\\\",2):f(\\\"\\\"{biSy/QvTw>aQChbi>vb5*Bx\\\"\\\",2):f(\\\"\\\"{b.T\\\"\\\",2):f(\\\"\\\"{:K.tb;=L<LNhbet?NO8\\\"\\\",2):f(\\\"\\\"}=evZaQaW9bbTaT7ep4\\\"\\\",2):f(\\\"\\\"}-pOHDTzbWaZaM|Q6H4Ga<Fwuoxt+g8s0yu9K7p8HhbNadbqqSCA,O|>=gbfzSaX>SYw\\\"\\\",2):f(\\\"\\\"{UnA75,Na,KTabbr>jsx5mDAaUnA7cyf6a\\\"\\\",2):f(\\\"\\\"}a4bn:6blbe<fwdbc\\\"\\\",2):f(\\\"\\\"{@Blrtb;4HIFI&6c^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'dIIPal>cbh5SXu8Pv8v8Wt.Y;y?\\\"\\\",2):f(\\\"\\\"}>Fa1x:stEx8RRmtO"));
$write("%s",("01wmOzg.0\\\"\\\",2):f(\\\"\\\"{/Fp5by?6bzLhb@a\\\"\\\",2):f(\\\"\\\"{b\\\"\\\",2):f(\\\"\\\"{*vb;0Uyl121i>f3HE@Ymb4*M\\\"\\\",2):f(\\\"\\\"{At<;F<jZabJC-VJC/bky\\\"\\\",2):f(\\\"\\\"{.ab,LCatJ*bl17b=abbo|Z=o79b1KwbN;RaM\\\"\\\",2):f(\\\"\\\"{OX8l,bFaqxOGqx-bE\\\"\\\",2):f(\\\"\\\"}>ajJc,?a@>7b=p1=/ydO\\\"\\\",2):f(\\\"\\\"{b\\\"\\\",2):f(\\\"\\\"}g4Yzj6r:M=L-b?2s1*Cl+Qa*b*bRwQqB?hbCLh/|5u5ebSsd7cNCtmdK7YadD8bYHQXG\\\"\\\",2):f(\\\"\\\"{duRwh/q+-n\\\"\\\",2):f(\\\"\\\"{/RaEalb;zSpty.bYH.0lLJdwaRa/lYamLOa2,\\\"\\\",2):f(\\\"\\\"}bhb/iVa/q53afdfb-b>pZaJ4nWkbPwCr74-LZBmL+DQaC3Pa7..8Itiy/bZa0bRDC3Pa@A<5C|>aGS=aKEyDab0wN5kb?-6zUa=a=aUaCIhb+cfbcNG-*==a;KZ\\\"\\\",2):f(\\\"\\\"}XaQRe:;@hb4Ai/gz@a1L7>|2c3@agqT/Rw|H=\\\"\\\",2):f(\\\"\\\"{dJ4smOtFbS@1k-bd8s=\\\"\\\",2):f(\\\"\\\"{Z5cbgHdDkbyBQao5qRcJOl13s49KB4Pak-x-RkQaM\\\"\\\",2):f(\\\"\\\"}fs+Tw>d-xbTacbyHEs4Ye<VPh7tv\\\"\\\",2):f(\\\"\\\"{@GX4"));
$write("%s",("byrUtKsN\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}=>8w?iueM|\\\"\\\",2):f(\\\"\\\"{CB;Ud^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'bD+bwbiS5bSG5LDLHw-Lfp*bgzCa2bF</nQaOax5Ya@\\\"\\\",2):f(\\\"\\\"{wbTa-s.QgWBBHw7q+Tlb9xSs:TOWK:3p;r7H51@tcJ3IRk\\\"\\\",2):f(\\\"\\\"{bD\\\"\\\",2):f(\\\"\\\"{,K|D1Y?aPugrA-tbF-:rWa;,Au>7q3cNbFH8m8<wbFa>=/q04M:oi7ueMn|y-e9z+3GkSfwdbqx7bUzu\\\"\\\",2):f(\\\"\\\"{Xa1KffKhzb|b8<qu*E>a,bmb-iQagPRpX*r2Va+6/b62vWOMb\\\"\\\",2):f(\\\"\\\"},RRt4wgZ*bZas\\\"\\\",2):f(\\\"\\\"{fxJwEaHGZ\\\"\\\",2):f(\\\"\\\"{xTWaOa\\\"\\\",2):f(\\\"\\\"{b4G\\\"\\\",2):f(\\\"\\\"{/m-\\\"\\\",2):f(\\\"\\\"}bhbKv\\\"\\\",2):f(\\\"\\\"{/m-+r1bgOnu*:5weA(6cCavbQaOaf\\\"\\\",2):f(\\\"\\\"}i\\\"\\\""));
$write("%s",(",2):f(\\\"\\\"}hbny1-3ys?q?\\\"\\\",2):f(\\\"\\\"}5Pw<z,bCLesab,1y;6JJzmbZa@x?aUazvm-\\\"\\\",2):f(\\\"\\\"}bVab4a;cpW1bgO++Da\\\"\\\",2):f(\\\"\\\"{bywYa-b?aJq<ruhrU\\\"\\\",2):f(\\\"\\\"{bhpsy2vPv8vRatbibN,BzZaf\\\"\\\",2):f(\\\"\\\"}1b3\\\"\\\",2):f(\\\"\\\"{1wZt6zJJlb<zA3<zf\\\"\\\",2):f(\\\"\\\"}1bKRxbn|St2DHGhba3<-R3yb++I+<wjTQj;:vb4w2wK2jBsPl14wdI7\\\"\\\",2):f(\\\"\\\"{|b*wbb6blOEy/9G5lb\\\"\\\",2):f(\\\"\\\"{32rAJ,K,w4,mv6H\\\"\\\",2):f(\\\"\\\"}w1\\\"\\\",2):f(\\\"\\\"}Crp54wVfouf\\\"\\\",2):f(\\\"\\\"}Ywn2\\\"\\\",2):f(\\\"\\\"}g\\\"\\\",2):f(\\\"\\\"{bo|QavfXx6b\\\"\\\",2):f(\\\"\\\"{b1b9x0-FapkhbRaA|WSczZas\\\"\\\",2):f(\\\"\\\"{9\\\"\\\",2):f(\\\"\\\"}P@c|buqpka>4tl2FwCr,pz1sM,wJw\\\"\\\",2):f(\\\"\\\"}w-bQZlb3bovky8wSaGw\\\"\\\",2):f(\\\"\\\"}gybgrA->8Na<ASrBplpNa\\\"\\\",2):f(\\\"\\\"{b<58bBBVImbb*AA/qtvV5NalBbnjbPN1x*sSu>q:@xvGaJEi3aacBvSwR72bGiN;5W4bKXnztbJ9PaAa|bCz>abb8s+6hGNvybh=6-gv0.h>hG@aq.Cr="));
$write("%s",("ydon\\\"\\\",2):f(\\\"\\\"{:2jEQVUxAak5QC@;m6Pan\\\"\\\",2):f(\\\"\\\"{h;atWas<P.tb7Ig8+bR5w<xwF,Ba5bS6/b5+NaH9LuabiGbb3t2\\\"\\\",2):f(\\\"\\\"}=phb6*\\\"\\\",2):f(\\\"\\\"{bfbup\\\"\\\",2):f(\\\"\\\"{bHj1wZpTOZu-VM\\\"\\\",2):f(\\\"\\\"{Za,6czb\\\"\\\",2):f(\\\"\\\"{WtEtc/Ok,mE.>z=K=mIM=3tJ=IxcLR9O=ybfb+lVa|=nxVa4DmbZA6qfbw*arC:6z6pS6fCYZYab=UaWai\\\"\\\",2):f(\\\"\\\"{RaetZBIrA9T-ybfb3bF=|bk^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fla\\\"\\\",2):f(\\\"\\\"})36(f\\\"\\\",2):f(\\\"\\\"{#,43z3m|a7693(f\\\"\\\",2):f(\\\"\\\"{#(ntnirpn\\\"\\\",2):f(\\\"\\\"})8402(f\\\"\\\",2):f(\\\"\\\"{#)K34SbKM\\\"\\\",2):f(\\\"\\\"{fbFaRROXTa-b9bub7Ab-/8M+B?Fa<DdrGaJS8b1K-WGX60fbt+>atF:KOXZpzvyKYHj\\\"\\\",2):f(\\\"\\\"}Hu>aGX80ffju+vt|\\\"\\\",2):f(\\\"\\\"{bSpPaQaS;ILkblDYahsRamtokOG:h3=XaA+Jd4bSc7b4=EA50Cr.bNaJwk;HrCaNRb\\\"\\\",2):f(\\\"\\\"}tk7b=aN"));
$write("%s",("2M;hYgfa\\\"\\\",2):f(\\\"\\\"{bM.5BEd[aCa*\\\"\\\",2):f(\\\"\\\"{nut6;y>aUzVa?aozSaK<+x|bIuRaE@p>E@,5O>/b;Huuyb|bIuM...Y@rOd8B\\\"\\\",2):f(\\\"\\\"{Z@T=@6<DW2fbGNRaPwu-M3avb>@S7Hrybqql>;1mbUaWa7bS.4mGaXCvblZd@X>E@lb;3JAy2gA\\\"\\\",2):f(\\\"\\\"{Q/u1jtbs2rzUzVaP-H-WMU.EaSambK2OadHM\\\"\\\",2):f(\\\"\\\"}PMGZX>Z@7t6ipU8->aiDz4aQa3bl>xpTau03b82\\\"\\\",2):f(\\\"\\\"{P-.0@x@Y,|=@a*xIL5b@;V<2A>63yi;QtFAEaPaL@Ru1/nF=p0YdbrACjnjIR|6c|dSBA\\\"\\\",2):f(\\\"\\\"}Pa/bINIq6puptkZapRwbSBKR-sRpQV1-UagDrCg0QZ\\\"\\\",2):f(\\\"\\\"}g>kw/TIiy\\\"\\\",2):f(\\\"\\\"{YlNrCfr+bZa0piZ5+tCgwPGVyg*Rqwb,beARaEaPa+bDa\\\"\\\",2):f(\\\"\\\"}8fbwbj1\\\"\\\",2):f(\\\"\\\"{Ie7vb3hJ.w>1bIrETIrb*7IvbdF562P\\\"\\\",2):f(\\\"\\\"}vkby9<D\\\"\\\",2):f(\\\"\\\"{TrsCyDy|9<<\\\"\\\",2):f(\\\"\\\"{jhbN5SWgb\\\"\\\",2):f(\\\"\\\"{RPBccksl>X*5Lju+vYa50CrR6aqXpo4?a,dCrJr57b\\\"\\\",2):f(\\\"\\\"}ab2\\\"\\\",2):f(\\\"\\\"}5bPa"));
$write("%s",("\\\"\\\",2):f(\\\"\\\"}=WaV6z:\\\"\\\",2):f(\\\"\\\"}/Es\\\"\\\",2):f(\\\"\\\"}/Nag/?Zdu7wMtWaC/K.Zo|=Es\\\"\\\",2):f(\\\"\\\"}/KhWa9ymb\\\"\\\",2):f(\\\"\\\"}u/b7-Zaz.2+>k3>&6c*dVatb\\\"\\\",2):f(\\\"\\\"}5|9zrBpUv:-\\\"\\\",2):f(\\\"\\\"{T6bg*WSnqWSIr6hWab9GZ;7@a4*TaJqiyS.s++dmb2Doxi=K+ubJ.Wa9yAsvM9bB3krQv1bvC+TB:H\\\"\\\",2):f(\\\"\\\"{Ya\\\"\\\",2):f(\\\"\\\"}wY*1*9r82h2kGyX55pGb6++vM\\\"\\\",2):f(\\\"\\\"}bTabbxs+6hbBaAJmb6/=BEp2-Ua1y53gvt4-b\\\"\\\",2):f(\\\"\\\"}zJQDaV5>aWS7bb:\\\"\\\",2):f(\\\"\\\"{b+;7w6b-.7btIPa:t0IF7=M.b-V*\\\"\\\",2):f(\\\"\\\"}QDCrq|7t5t3ts\\\"\\\",2):f(\\\"\\\"}wI5bH*<HN+*;6z6pC3Wa?ad7lbhbNajbNXYaCa6HmbK9130bG|Aa4Ehw=pf;q|etYatbZ8Kvkb1w06ccafbWTega5D>6/nh<aKaRhRajrX>R+/OUi:5Gv4wkb++fbRiWadbcbc3hwc;dbT7ubV*v=\\\"\\\",2):f(\\\"\\\"}Tzjt8<9hb9xCC\\\"\\\",2):f(\\\"\\\"{bQtUXI3cNbiK>aPa1bvb-retRkt0nW:qZa3b-6XaPN5wA-0qRphbMxB1P\\\"\\\",2):f(\\\"\\\"}eNs?q\\\"\\\",2):f"));
$write("%s",("(\\\"\\\"{m25bMS<sCs?S6J4betlvIry.Av0E9=jTibX+9fH0MPhbx\\\"\\\",2):f(\\\"\\\"}9yKv;PdbFan1y5cbh6=aC\\\"\\\",2):f(\\\"\\\"}Ta7bY@KvPwy5cbkTovBJcW;7dbCaDaKvjbq*+>C3cuajbwb\\\"\\\",2):f(\\\"\\\"}vBpUva@4wUi9Z\\\"\\\",2):f(\\\"\\\"{0(6c?gUvld\\\"\\\",2):f(\\\"\\\"}w1K<vjb/1jK6bFat5hbA*dbDu.M,M+vOXTaNJwA0>m=mbn=t0n4jsK92@y;Ya\\\"\\\",2):f(\\\"\\\"}+>aoJ@P0b6t=al>9,,bj\\\"\\\",2):f(\\\"\\\"}Va\\\"\\\",2):f(\\\"\\\"}+/HpF?<Ea?rr5\\\"\\\",2):f(\\\"\\\"}H5,RaBp6p6|4|*\\\"\\\",2):f(\\\"\\\"}Is*\\\"\\\",2):f(\\\"\\\"{9uRa2TeThbDn4bo\\\"\\\",2):f(\\\"\\\"}:22T-KK@-sCr/b?1M-futw:3Wa?IXp>RhbBaZ<9s\\\"\\\",2):f(\\\"\\\"{@+0TJs-Oadod7Ga:8ib7Io\\\"\\\",2):f(\\\"\\\"}dbdH.zVj1jVaRkQYmIwyoyDnS6-WWaQRcGMx-40I*J/Hrz||Y@X,GA1yG|wIoIN02bmbDaZa/uI-DaLM1Cy4uY:SabU2.8NrEFSc+6;AR|.dlNxbQ>puEF=>mDPw;pgwK2CafwfbCaJ/XYab.b*\\\"\\\",2):f(\\\"\\\"{lb76R|OhCaEFxbE-j-cbS;d/nW8blbubSaZF0pD<ybVzab.bVzw5asOvQ39rf"));
$write("%s",("bN<YaNrbR6soyZ\\\"\\\",2):f(\\\"\\\"}9qNrKONr\\\"\\\",2):f(\\\"\\\"{bZ:8hz:2P\\\"\\\",2):f(\\\"\\\"}vlb+bBa=|EFxb6uer9qNrSasq,KUavs@adwywfbh7;p:r;pGDK.H3SadpCakbPa3pQvhbJx01P\\\"\\\",2):f(\\\"\\\"{B4OlW,v=K7HJ\\\"\\\",2):f(\\\"\\\"{bBJA-<6?aB1DaW,v|/+Oqk\\\"\\\",2):f(\\\"\\\"}ubhMfM@aabR+fbFaub>McME9cga\\\"\\\",2):f(\\\"\\\"{bPacMe3aEac8F,:qYA2w972bOab-pxN02b254pt@I00bo12w;:SaecD7:pryuZhbEa:ffp.7jK8Hcycwzt|ebbqF\\\"\\\",2):f(\\\"\\\"}9;Ra3tmIE\\\"\\\",2):f(\\\"\\\"}*sy.k\\\"\\\",2):f(\\\"\\\"}ebZtVvRaCBAaSzETy<WM0XP-2b/bk5n?+T4tHI?acbj:Fa8sH\\\"\\\",2):f(\\\"\\\"{NGo|yrIS9A:Y1y=t@\\\"\\\",2):f(\\\"\\\"{Ra71\\\"\\\",2):f(\\\"\\\"{b,xQvrNpNm2qxUaUXg4?acb?aqClb,3g|X*EA9bsLfb3bO=|bZaSTRs3=diyby1mxaw@57,g8jb20.ThbJ76b.w:sxr8bZaebibB4afaiHPvYQ9d\\\"\\\",2):f(\\\"\\\"}dnt2rH-I@+s6-Va<=ynPaJ4;pVaMQ0*xb3=2W6iITwb.;zbfuYaNAO?nY6btE>a|wL|91bd0bXtXatyk+=|814>39dbdHbOvz7t5taZX0"));
$write("%s",("Zsoy?a>|4|6bcbiS+sN<b>Tayp2PEas@aqh-,bputbDa0bO>h8mN-KWaW.+tybybBa3trRE|*\\\"\\\",2):f(\\\"\\\"{1Kp5mt/b;Y5b2r=x4UYEbqlDD4Q39=?aCBfS>ABapGtlMp7AhwPv\\\"\\\",2):f(\\\"\\\"}bVa.\\\"\\\",2):f(\\\"\\\"}vxBsB*;X:-NXtrX>.b8CK7WMh,hbeyCa?abbL0\\\"\\\",2):f(\\\"\\\"{rGjmbbO3ygD4bv|Nd4b.;xbNa9,9T0v4SLT2w4w1bO=c?RFREIr5bH8*pTp\\\"\\\",2):f(\\\"\\\"}w:qL;Q|FAf;h86bw@ukEaPaSiYa+bLLRCtU8q:PV79>yb91*b<z|vnvDDJz5p|\\\"\\\",2):f(\\\"\\\"}6-s<bbTauhrUhz7-6/B*xbRCtUubZa;3cmaC|VYkbxu6b8b%3a^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'bOXPvYamdNa;|tUFy:PV7Ru/wg\\\"\\\",2):f(\\\"\\\"{T\\\"\\\",2):f(\\\"\\\"{i2.ubbTaj2h2NXCr>>ebdx8bJ7-M\\\"\\\",2):f(\\\"\\\"}b-bgUbJ5\\\"\\\","));
$write("%s",("2):f(\\\"\\\"}zA>Ru5ebaxbqwb>s.bT=,rxwNqdW<O3bfsQts0hbCaeqUnEBbbT;.r.^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'GdY2y>Pw:Gf\\\"\\\",2):f(\\\"\\\"}CaBWcy6bCay>WZLP7qSZTa7wvbts\\\"\\\",2):f(\\\"\\\"}gc8h2HZNagb6i8?y++\\\"\\\",2):f(\\\"\\\"}CCxbuvU2*b:M>==Det4s8b7sdbtvs13+F:w>fbgbr*K7o|3D2Ns0M7rshbZa?y3L.qebML*My<lb9\\\"\\\",2):f(\\\"\\\"}jr-vYE0bw*>yMLuxV77<fb@PdbcL4=bb2qVaYH.r9b\\\"\\\",2):f(\\\"\\\"{bAu876zGasG+b<z;<A\\\"\\\",2):f(\\\"\\\"{y.p0+bJY859|l6ewgcpFyMbbR7BhVyX0RpX96iL+=L9KVuc4*bBaAawv+1gwMC.bSw5bdbaK9LfbYa|bxboz13Ga,9S=TtOyDOMKb2|Wu..pSL-b\\\"\\\",2):f(\\\"\\\"{*Htu=\\\"\\\",2):f(\\\"\\\"}b0.h5wrdr9bOW:2fjr\\\"\\\",2):f(\\\"\\\"}qRYaWuju@.y\\"));
$write("%s",("\"\\\",2):f(\\\"\\\"}G3vb.;13STebcNgbgb2bTaNa:Ehu4Fkb9b?sV6DDyv>aRkJC;0BpYa=aUi1jRi>a6i:0@rGaTVCsB9=r>ayV9bxb=JICeX+lIkxucW\\\"\\\",2):f(\\\"\\\"{rhuFuBC.bD:A1H1kS@0p>TpNVtrY5b:br+FVAqvgbdbD=|vNxSL+bCa7bNV6b|2gb-bEaybi9Fas0Nwp0yb3IH:2+guiS.bdb->oHur2bk5gb-wQ|pyhwXSV7q|Bvab-b=s;sKr=a-b/k5C;S7UXapiOrsW:Kib=at4|b||PhXatbfbFx,bI0hbP:Pa\\\"\\\",2):f(\\\"\\\"{b=AFjctub-V+@J-GEOap/2+s/eL,v2NXaEsJiE+:r.ptr3mdrE+SLDAib=u1xy96iTC7:0*Hkp-UaINLir9O0m6gxZr8*hw=udVp/XIXaSagwBvd|ky03SPYS|f+E6Flq@0*7ok</LLctn17>JC4*K9ySfbs4UtTyYEx89b3+\\\"\\\",2):f(\\\"\\\"{bK9kb?/Dpus3sR7mslNtE6+=zl0,b8+z>D2Oa3IiQ*:551jhUaPPEFD9bgb=RTaE+>-LM?QC|@aYNYqup9b@r*bHIb1wr0b?2YRnFg*Wat52jlD\\\"\\\",2):f(\\\"\\\"}b7whbG+w-\\\"\\\",2):f(\\\"\\\"{uCr0TaSUa8..xE-fr?rbb@+FI<sH*dt|bj\\\"\\\",2):f(\\\"\\\"{Bwfbv=fKnq<P|bcQxwl|w?8<3bZa:MCrH1ATO>kbYa*b0S1xm"));
$write("%s",("3p5Qv5+B7D,KLkBEaQv-bq/-G.TmLTaYwzbAaebwO1,,b<\\\"\\\",2):f(\\\"\\\"}2*TaCr5+zNzgwIMCh|OaQtA*e4dbOaE.gxMuub6b@w?a,COq\\\"\\\",2):f(\\\"\\\"}b5ww,iSFSASEagb6bOaE+GD1bIN*rQa:rh|Uaf:6izuOa<u4bMuNGlb6ik>hC6/5bLM|?-ACOIMxrWrl|\\\"\\\",2):f(\\\"\\\"{Qzbibkb>0c:gsWB>0B:OqDpyjUaY5=4Lofb;zyb<vzp8=@>6bh6Ea3\\\"\\\",2):f(\\\"\\\"{rG2qB--bB:FaG|/bA9FaWaZK,bebeN3bn2LuF7/bBzbsBa3bGr9br>\\\"\\\",2):f(\\\"\\\"}7N;cb\\\"\\\",2):f(\\\"\\\"{zJ2QCYH<;s.AAy?aPTODaebFafbTQ.2QaGsq,yBo7g//p-O+rtx24h,R5iB7bLv2Q/--sab@0s4cyzb=aNx5mv+*\\\"\\\",2):f(\\\"\\\"{?a0b*\\\"\\\",2):f(\\\"\\\"{Z;wbNajpTqRqPqNqLqqu@9s\\\"\\\",2):f(\\\"\\\"{Ba*b8Qtb,54bZ:d+Da|bi8L;xAJ,EaBax8v6Caf|0-,z;KyI+Nd2MII6?GLMhw6?lErqD4qF*b\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}-Fqvaq\\\"\\\",2):f(\\\"\\\"}Cbb\\\"\\\",2):f(\\\"\\\"{x?6*D1bibC9KEu2PaTa\\\"\\\",2):f(\\\"\\\"{bIpGpupl><7SOkbValP:uek;-x\\\"\\\",2):f(\\\"\\\"}Urvb3Iyb"));
$write("%s",("/Obbgx=uyrw>e3O=yv@,HGNa.d1b@D8bgb=u/q=a?vaxCakyN+-vOagc.,k@G,Nwo7abk3hbNqe,Xac,mb3bI4Q8yn7;e:+1BqwbyMM.e;1Kybm=exi/fEO>6bybjbs,as6uLDx?Faf.k5drd8k@<a,1S0PavFn37vy,pi7,W1,,kbD4MsXaVaF/+*kb<a\\\"\\\",2):f(\\\"\\\"}xmDo9Fsjb?4WaYaEad2E6AEH6o;r;IKJy.O+6eih803ubh\\\"\\\",2):f(\\\"\\\"{jrMw1y?40x1b|bYaw*oA,b\\\"\\\",2):f(\\\"\\\"{bFaabzb>ykC=aQxBuk:-64u8b<;iK:;8;s</<R|=1Bv\\\"\\\",2):f(\\\"\\\"{bCaJ9d.\\\"\\\",2):f(\\\"\\\"}v|*@a>-p2kbjbTambC7VaBDl/qHaL0u.uX<mb6bh/*.C,NqZ<lbdbD,.u=NV.S9J|6-9=|=.bg07b5xcb3bIk>F?1avMxD1R6abZ:Q\\\"\\\",2):f(\\\"\\\"}gDs\\\"\\\",2):f(\\\"\\\"{BsG-p6EHy7hb87PafILBX2T-Ku9\\\"\\\",2):f(\\\"\\\"}L4jbabf|tbR7TlRaKuT-H*5zm.+1+bxuabA|h,tEX6X43bozOaawp3uzPaNaB\\\"\\\",2):f(\\\"\\\"}6-4aJM\\\"\\\",2):f(\\\"\\\"{4JI@aRD16X<Gx9f<0<aEaq+7.Pabbfj?,bbWagw*j5Kub6u\\\"\\\",2):f(\\\"\\\"{+OafLdb>><>\\\"\\\",2):f(\\\"\\\"}b:>@+wb*0@;tv,7Daz=r"));
$write("%s",("\\\"\\\",2):f(\\\"\\\"}tbP\\\"\\\",2):f(\\\"\\\"{ML2bD\\\"\\\",2):f(\\\"\\\"{Oa<7dH?se30bjAk\\\"\\\",2):f(\\\"\\\"}1y>8>aIL.bjAyb3bzvcw8rfu0bg9k+lrvbE+z\\\"\\\",2):f(\\\"\\\"{OqE@@F8bwbGam|5b8Lz.2v:rjbbbQ\\\"\\\",2):f(\\\"\\\"{@FupzrVa\\\"\\\",2):f(\\\"\\\"}bp0mLzva?+6s+N4\\\"\\\",2):f(\\\"\\\"{bIuNa5tYaCrC79z\\\"\\\",2):f(\\\"\\\"{b2bS+6baxBh6*gbi|/E=afbk\\\"\\\",2):f(\\\"\\\"}c>8bUtubcwUaBh4b<5R9p6Hxk,UAX>vbPv8b<a=aQa41\\\"\\\",2):f(\\\"\\\"}bCx/-9Ko:m:fb\\\"\\\",2):f(\\\"\\\"}bquotJK,-p;,|d2LIuc42*zNq;HbrBujJ4|H\\\"\\\",2):f(\\\"\\\"}S3xwuA0bZavb;3FaIyPs<s4b?-+byH/qQz7bzb1j,b3DNCH1mz\\\"\\\",2):f(\\\"\\\"{.Ar=-s\\\"\\\",2):f(\\\"\\\"{;pWhcxubtE/HVHyn?JwHvbjs\\\"\\\",2):f(\\\"\\\"}bAIR=Fa=7B\\\"\\\",2):f(\\\"\\\"}E.YaYa@a2De9lHfC4=FaTaUa5bnz\\\"\\\",2):f(\\\"\\\"}b,bOidbbr9b<au-g*A\\\"\\\",2):f(\\\"\\\"{u.0E58?aFaT|R|hrVaVIoJLu5+*y\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"Y-eb4zO>T=Xa>\\\"\\\",2):f(\\\"\\\"}@a\\\"\\\",2):f(\\\"\\\"}l|r5wn.5n"));
$write("%s",("\\\"\\\",2):f(\\\"\\\"}bRqCa+b;wxz9zfwmz8-Sas\\\"\\\",2):f(\\\"\\\"{Va\\\"\\\",2):f(\\\"\\\"}H\\\"\\\",2):f(\\\"\\\"{bq+hb+6-s*5.bs\\\"\\\",2):f(\\\"\\\"{Ra*5H0AINa8b8bCaEp1b|rmD@a+l@aG.Oavb/p|hOy--r=O/=Gdb-bBadb5EBB\\\"\\\",2):f(\\\"\\\"}b1jybbsFaBztImbi.WB|bn=Eamz0.ei0bQa.bFag/Oamx\\\"\\\",2):f(\\\"\\\"}8hI1bW\\\"\\\",2):f(\\\"\\\"}yAT3dbSar*Fa0ljb.b*bgray?s2b=7>aRaF76iUH+HH\\\"\\\",2):f(\\\"\\\"}7bmqRaPaTu4|W6cb0HgH\\\"\\\",2):f(\\\"\\\"}8Fa+GV-+H6ss.abwHUfBabrVn0z0lhH<aSa5b=:6llbs-IrdrNqUaVaZaBBSaeb,bn<l/D.L,Os>a\\\"\\\",2):f(\\\"\\\"{b,yjbk@Zo.9Vaub\\\"\\\",2):f(\\\"\\\"}p02ZaSaA|xb?aS6=aF75bW,<7EAxbUaZ=1bAa\\\"\\\",2):f(\\\"\\\"{bybzbl/4b<a>sAv/bM|ypBCzb>a6FRa=pb9-bFa2bdbQv|bS6Qa6b@a5z5bKid2,?4CJm?E/k=E;rw>ZaDpejb\\\"\\\",2):f(\\\"\\\"}YFMr4w6ba7+@j\\\"\\\",2):f(\\\"\\\"}9\\\"\\\",2):f(\\\"\\\"}Za|\\\"\\\",2):f(\\\"\\\"}qpab@\\\"\\\",2):f(\\\"\\\"{1w>4n6Na>=d-up;|m3jtE<1w4vjb8FL;-bUz\\\"\\\",2)"));
$write("%s",(":f(\\\"\\\"}bw58bebKqgwou42ib45=aEa\\\"\\\",2):f(\\\"\\\"{bQ9O96iM97bK9IjH91b>a4e<ao7LDn<L|z*gbL-Psrq?aX2-blbf,+u6i5:mq<hbbfbP.2b\\\"\\\",2):f(\\\"\\\"}=4bPBAA9bCBxus+Fa220*YAO=on*v\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}v+/s?6wb42ubO:gDUa7b\\\"\\\",2):f(\\\"\\\"{@|bbpCrVt8qDE4b\\\"\\\",2):f(\\\"\\\"}=wvwD@an:BtH9;1|b7,jbR|21p2d1gD2DBazgoxBt=/6ihyg:Ga8:v+x\\\"\\\",2):f(\\\"\\\"{ibOyZ1+?1k2CBi0CFaZBh,u\\\"\\\",2):f(\\\"\\\"{>aYa|5y9tb<a<a>alb\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{0v=,+1*bwbzsKDp2gE=>ebPaM1.9tbD<cyXa+bBu3j6btbV;3bEa/<>aa\\\"\\\",2):f(\\\"\\\"}hr0vI+x*ybWaG\\\"\\\",2):f(\\\"\\\"{e?Zs=wtqevUa>a\\\"\\\",2):f(\\\"\\\"}bCa<ayr=\\\"\\\",2):f(\\\"\\\"{QaQaf:wbC|db.b/D7bo:Ca=t3bb:y9fbabBae;dkA7ms0b3:tu\\\"\\\",2):f(\\\"\\\"{bAa0-D,3x7:K@H.28Ca|2db87l>zb:pvb-6K9DyQalbxb+lu.B7Qa4bVxTxUa1bkbf?aD5b>aUaZa@B6i0<J9F-Cr5babNa/b<ap5-b6bjbVylbXA995+acp0Uyu-.b?sm97qQ3"));
$write("%s",("vbu-dsm-K+UaC\\\"\\\",2):f(\\\"\\\"{Bi+4,A<m*A6k|A81Vy6bvbFa0b2bo4Zp\\\"\\\",2):f(\\\"\\\"}gK+64:31bJw4uP\\\"\\\",2):f(\\\"\\\"{@a?ad|7\\\"\\\",2):f(\\\"\\\"{M3RB+b\\\"\\\",2):f(\\\"\\\"}bo5VsOaW6ebKfPq?s+1WaUa/+1wibzbJ|.b1bBa1bZaLsm=Xykb5b*serruTv:pgbxb.bTa5bfb2@yj\\\"\\\",2):f(\\\"\\\"{bu+Y@x\\\"\\\",2):f(\\\"\\\"}Fim-Pa<a7>|h2v87A9z>|x-0>s5bS7?19=f-nuq|Za\\\"\\\",2):f(\\\"\\\"}gwp2\\\"\\\",2):f(\\\"\\\"}N9Y,m=Huy.NrJw+z2u6i\\\"\\\",2):f(\\\"\\\"}m\\\"\\\",2):f(\\\"\\\"{babf:K0S>g:/r@aJzjui;ybOai;*bVx?uvbAsUfr?QaxbmbL0G.Nq@9;41bhbSaQaB\\\"\\\",2):f(\\\"\\\"}R7/bvbUnjb0bzb+b9zNaLpWacY2,jb\\\"\\\",2):f(\\\"\\\"}bO+AaD5MtvbOy\\\"\\\",2):f(\\\"\\\"}-q;9k\\\"\\\",2):f(\\\"\\\"}?H6\\\"\\\",2):f(\\\"\\\"{?=-L;ab2bibz2AaM,nA8bdb=t2?bbVx2@FjYaY.5/t\\\"\\\",2):f(\\\"\\\"}.p+bG=JzUid+P@@a+bV*b5.uT<i1@@F-+xepX>6-@aVa3bzbCrWa8bEaNq?aw@|7E\\\"\\\",2):f(\\\"\\\"}d/bbubD5=pxb*bP:H*@aN+Ea/bWazbBzEwUzM.M05b+:,zx"));
$write("%s",("vabSxi>\\\"\\\",2):f(\\\"\\\"}6Tz\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{.d4bBag<6iErcpp65xxrebz+Jzf@D|2jwb914;eb3bmbN4Q\\\"\\\",2):f(\\\"\\\"}<aZs4t5|Vz0w9b-bXaS;M-n<*xR7l/;4er**q7cbX*fb?aR|g+:qUt6b0vq|pswbapWtK0.9s:4b\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{Nv,bAuOyQ/*46kG6d2p=Jxtbd1xr\\\"\\\",2):f(\\\"\\\"{bCrK7cb.bH\\\"\\\",2):f(\\\"\\\"{.be:A|dbZ8x8.wg|cxG>=a85abL9Gv6bT;V>CrB4xbL0DyI0+bab7|>azsRrt>YaXaBqr6Tat1q7k:W4Y=SqkbEu6s3b@.Q\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{yAaD2ub+vx8abAag,J,sqNwibcbB1Ca8b,bJ/;rlbSr>=kbUqC9TxS=gb/bRaG+z3ubCrQaIqgb+bG.|s0bT/vbZacb6bQayjE.o6Jw9bZaNaVa4bCaAapuCaek<7Jw5bub3/Fax2BpX.8bj\\\"\\\",2):f(\\\"\\\"}-7.bL<5bBa@aUaRaoxU<Aa3bkbqq.b\\\"\\\",2):f(\\\"\\\"{:OaV<Bs-.6-V.WaSa\\\"\\\",2):f(\\\"\\\"}/?aT7K.Irkb2rd2J6x4V8n;=x|bRa2j:rK.Aagk3sn4Rs=/R3BzK2mb94Ea?9Ta@aUzK2P;u5PhQsmbv5PaWa-.cpCsY\\\"\\\",2):f(\\\"\\\"}Cr3bwb"));
$write("%s",("nrt1Kvb<+basEpvb<ah/@;0bEa,buxn*l*\\\"\\\",2):f(\\\"\\\"{<ZzlbkbBau.ds|bvrH9|bkbu8wb\\\"\\\",2):f(\\\"\\\"}:C;2zmrr9gbnv7bg:b*0b*bJ.Gjex\\\"\\\",2):f(\\\"\\\"{u07ub0bPasiP-AaUa\\\"\\\",2):f(\\\"\\\"{b5bCzAt*bZ|N2Sat9;p@aqqPaZaub|bVagz4;1/h2k\\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"{L4Wz?rRaDo4u;1Xaw+1yNaEa6b/xib9babpvY,L7nrkb;*@xUavbQ\\\"\\\",2):f(\\\"\\\"}j1w|b-ebQsZ8PaYaz+|oH6c2\\\"\\\",2):f(\\\"\\\"}4a2W8Jztb8b\\\"\\\",2):f(\\\"\\\"}+Zalb|b4bcbtkUax8\\\"\\\",2):f(\\\"\\\"{vcb@+,bDaTf<84bd|\\\"\\\",2):f(\\\"\\\"}lDpFa/b2.dbdbxb9bFaF|8+.bPrP\\\"\\\",2):f(\\\"\\\"}vbTa3\\\"\\\",2):f(\\\"\\\"{Nabd2wYasqybmb6iDt8bp2yupivuPv.5gc\\\"\\\",2):f(\\\"\\\"{rEa+*v*bb\\\"\\\",2):f(\\\"\\\"{bubUaEaebVa/p7bW.D|.x7bq.2\\\"\\\",2):f(\\\"\\\"}@aTaZa+bFqabwrNwH00bkbWa.02bDaIrgzi6SaWa2,/9am\\\"\\\",2):f(\\\"\\\"{bRa3pDa@zCr7rtqeb8bK+*bEx<7-bbpZakb|b\\\"\\\",2):f(\\\"\\\"{.WajbQ1.by+c3Dau9T/fbc8OaPax*\\\"\\\",2):f"));
$write("%s",("(\\\"\\\"}bZatbQan|h+Fau913Na.7Yjjb?\\\"\\\",2):f(\\\"\\\"{c35xl2abP0zbBhp\\\"\\\",2):f(\\\"\\\"{zb2+,blqTvyb1bv6mbV.dbTa/bVaq5Aamb|oT8F6e2D6Wa,uBag7@a<6LuGuUaubYu3bNp,bIu5bN|lr|7@s-8jb+8*b6i|8s-:hkbm8Na/8d1|bz6lq@abbtbwp\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{RaCrV,Vs4xD2lbyb/qgbKs1x/bfb51uv<a0bwoW,xpubtbTaE\\\"\\\",2):f(\\\"\\\"}z2-bubJ7p7.\\\"\\\",2):f(\\\"\\\"}m7k7b3ebXylbtbwbE7;1z,eizrQawbabar1rv|Ra5+8b3bXaibXy.pybhb,bUaq|wbwb?avbybiuoiEqgjebd1Cavb?ahb|\\\"\\\",2):f(\\\"\\\"}8b\\\"\\\",2):f(\\\"\\\"{b.pg4ubRaV,BaEywbY-s\\\"\\\",2):f(\\\"\\\"}xbY06buv=4Qazj9fBa/bEabr>a3bN4rsBa?t\\\"\\\",2):f(\\\"\\\"{xXalbWa,yib>ambCr<y06ab.6,6OyLyPyz4|4OyP*Y1*6>yDaubWatbfqUazbGpevCalbd\\\"\\\",2):f(\\\"\\\"{cbBufx<y.bn.71cu@aBaab=a3bopS01bE|Z\\\"\\\",2):f(\\\"\\\"}B.Pag,Aa/b>a+*9b2b>a5b/bCaA3Sa1b1x\\\"\\\",2):f(\\\"\\\"}lfbDa3b/bE\\\"\\\",2):f(\\\"\\\"}FaCrtiN+xb7b1b,dzbn1L|"));
$write("%s",("<yWayb9bwbIq\\\"\\\",2):f(\\\"\\\"{v>a*bybd-Ba2bj1|bub;4bbUzcb9rYaetCrQ1Jqwb0bWxZa-pBtD+7bg,jb=aTaeb-bVxmbcbAa@aWa=aSaS.cbebOaQaL*p/Rxbb9b621bD\\\"\\\",2):f(\\\"\\\"{9bNaI01hPaN3|wXaWambD4iyG-M3VyQagc4tubmbAa5b0bibBfl-i46b2bL,\\\"\\\",2):f(\\\"\\\"{bEa4bdb|bibS2\\\"\\\",2):f(\\\"\\\"}bQ2Va2ba.Cr=\\\"\\\",2):f(\\\"\\\"{r-ItBatb|bP\\\"\\\",2):f(\\\"\\\"{Q|db6kM/.|d2Ny5kN/Qy+-jceb1b7b,b6ix|ppeb.b738bzbOaM3w|ub6s/bBafb-,?,Rt9,4b*bT02b+bkbQa9b*0=|w\\\"\\\",2):f(\\\"\\\"}fb2r*bBfSaFabbepT0p3>aeb2bZxh2j\\\"\\\",2):f(\\\"\\\"}3eu+QaTaKqG,0b5|tbx2.n9,\\\"\\\",2):f(\\\"\\\"{b*bq3WhM\\\"\\\",2):f(\\\"\\\"{6bUagbBa32Cr1hZvFxybebz\\\"\\\",2):f(\\\"\\\"{M,LtXaGu7blpvbPa;|vbB2d/wp;1fbUa\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{0bubEaibtr>aybu-+b;-Wa*b.b6\\\"\\\",2):f(\\\"\\\"}pjlbexBhQazbcbXaTa4bq.abt1T0=/Rw4bg*vb:*7tlbevNaIj0bym?akbjz,b5bh.*bqpybdp0q3b>a?a*b;xxb\\\"\\\",2):f(\\\"\\"));
$write("%s",("\"}up2Na5xxb6bI\\\"\\\",2):f(\\\"\\\"}Cr*sXaFa4bus@.8bmbi1ot7kO*pw-|*-yqP/4t9171JxqvUq||PaUaxbbw4b5bp\\\"\\\",2):f(\\\"\\\"};zz1fbD*f,/bQaUqlbjbPa3b31-di1Sa2-*bab<aFa3bib:./bzrwb<a8uScXaeb0pk,V*q0Na*bRa.qLhyvNa0btq-qh\\\"\\\",2):f(\\\"\\\"{hb.bYalbz.Pa8b/-PqWa0v0bSaNwfp7\\\"\\\",2):f(\\\"\\\"{vbOazv?y0bdbgbWafbZa1bwbE\\\"\\\",2):f(\\\"\\\"}.bib,\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{bmbzrT+R+-q@0NzGaLz*sYaqqjbCr8b\\\"\\\",2):f(\\\"\\\"}05b,09bDav0,0.bz0+0\\\"\\\",2):f(\\\"\\\"}0*bDaW-@aEaW-zbDa.b2|Ea.b2qEaYawb2r?aOad,6/x/UaDnD-7urzOaF/e/a0D/B/C/=/D-ltcbCr>awbA\\\"\\\",2):f(\\\"\\\"}otT*L/mwS*wt|-qnlbM.F/@/\\\"\\\",2):f(\\\"\\\"}bR.?/Sag/Qzg/Qae//blb;-//ev5/8-1bRa4bzb0bRa/\\\"\\\",2):f(\\\"\\\"{Nq9b0bOrk\\\"\\\",2):f(\\\"\\\"}VaSad-ebEzZaabRas/3*q/6io/3bCrK.<aWalbRhL,Qa=ambfp=a+b?aSaQvFs3bDalbVa.bcsRa=a7bOaw.D-8bPhRa>aEaAaSa6b+b@a/pSaT\\\"\\\",2):f(\\\"\\\"{yb"));
$write("%s",("6-7.ynVzVtOs|*5bXa2sN+=aD-?a*.Sa>u@aSaAaWa.b9y:habtbAacvUu\\\"\\\",2):f(\\\"\\\"{pmbmbtbzp>a1bYa.b7bgv-b=a8q|bOa1b;|Carvdi5b8zRa.b\\\"\\\",2):f(\\\"\\\"}b\\\"\\\",2):f(\\\"\\\"{bynQa7uFapu+blp@xkbSadb0bbbSaTaOalbRa9bPaVacb-bAatbRaQaPa=aab8bWaejAaevtbBawbUaot+|qtowQ*/|R*gbTt?aCr2bSsNaxmfbNa*\\\"\\\",2):f(\\\"\\\"}|\\\"\\\",2):f(\\\"\\\"}h-?aPazbRa-b7wZaD\\\"\\\",2):f(\\\"\\\"{5bflebZajbm+0,VaFavbRa1y\\\"\\\",2):f(\\\"\\\"{bnqSap|.pix4bUalbib6b\\\"\\\",2):f(\\\"\\\"}ymbibCa.bOambOs=a1bUa5mEaNacbPhmbbpRaabxbEa0bUaFaCauv8b/b0v@aD*6s*bfbcbLxlbgk/bNq|v1bp+>a=xT+vuOaFaFagbXawbgbibdbgzjb3b@ftkPp5b<ahb-u9p3b\\\"\\\",2):f(\\\"\\\"{bVx1pWaEaCr+blbD\\\"\\\",2):f(\\\"\\\"{3bOl6in+lb-b=u@akbAaSwTa@w3+0**b>aOaAtkbOaWujbOa=\\\"\\\",2):f(\\\"\\\"{fr1hCa2\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{bUaEzXadb<a+bTa0v4|YagbabbbEsVabbts0bVa+bCr|rCrubkbVzwj8bwoW|N|\\\"\\\",2):f(\\\"\\"));
$write("%s",("\"}bSa0b-i*b|o/kvtN*MyrwRy*|8b@a0b>yA*Vaejj\\\"\\\",2):f(\\\"\\\"{-ikbr\\\"\\\",2):f(\\\"\\\"{+bvbI|lbmbDu1*2\\\"\\\",2):f(\\\"\\\"}7bqpeb,uvb/bCrVa0bOaXarqPa@zcp9bQaUxXa\\\"\\\",2):f(\\\"\\\"}b|b,bcbQa2\\\"\\\",2):f(\\\"\\\"}Z\\\"\\\",2):f(\\\"\\\"}wocuWaDaJxTa@yWa,d5baxDa\\\"\\\",2):f(\\\"\\\"{sDa6q\\\"\\\",2):f(\\\"\\\"{b4bfbQa8|7b=tZtAuCxIrQvD|7xOaxb4bxbybbthbPatbzbk\\\"\\\",2):f(\\\"\\\"}kbgbuf,bkbbbj\\\"\\\",2):f(\\\"\\\"{5bgbzbwpvbppFa?t?a5b|babzr*bsy6iprlbEadbzbdbUa|bvbAp-bOaCaR|5mbbbbNamb8bNa>a<ai\\\"\\\",2):f(\\\"\\\"}=aYa9tAubqhbWa?p6\\\"\\\",2):f(\\\"\\\"{zbXaXa|\\\"\\\",2):f(\\\"\\\"{bb3b<aRa6bBaeb|b7pTavbvbWapu<a1y7\\\"\\\",2):f(\\\"\\\"{0bvbwbtb\\\"\\\",2):f(\\\"\\\"{bUwAa>v1webzbfsmbbb,b6pQadb\\\"\\\",2):f(\\\"\\\"}babat?a@p|o6kutOystOyKy<axbC\\\"\\\",2):f(\\\"\\\"{@aps4bNawb9bhbfbjs4blbBa6iauUaCaWuEpZambSaY\\\"\\\",2):f(\\\"\\\"{Bahbzr5qtbNakb\\\"\\\",2):f(\\\"\\\"{rUqus,bip+25bNa-b<qMp8b"));
$write("%s",("OvOiVx|stbcb.vkbNa4bVaQa+bjbYjdbEuou6bKsOxcbIda\\\"\\\",2):f(\\\"\\\"{Pa2bAasq=aOao\\\"\\\",2):f(\\\"\\\"{JribSa8bOadbYyib8qxbAaNq8bFqSacbOa>a|b|blb1b8sEa.u4bRa\\\"\\\",2):f(\\\"\\\"}zhq+bVakbNzCrmbkvnj3bubPa@a9bRa8zhbyb6iHshzzb?ytsgbZa.bvz4bjb.qAaxjIj>afbibOvRakb2bBaubfbywEyVaYa2j6bnv3b7bdbabTa3bKqpy/bDa2bfbIsYaUaNv+bFaYaeb<y1yybAaXaab*bOa/b/b6bOrZa8b7bwp\\\"\\\",2):f(\\\"\\\"}bNafx1kxtkwptqwnwotrtjwub7bAt|yabibEa9f?y3tib3bYaqvmb+c\\\"\\\",2):f(\\\"\\\"}bDaiyjy,yRajs1boygb+y6idymr\\\"\\\",2):f(\\\"\\\"}bUn*bibev\\\"\\\",2):f(\\\"\\\"}bcrtb@a\\\"\\\",2):f(\\\"\\\"}b3bHu/bibRaUqSaub-u?sGaitSwCr\\\"\\\",2):f(\\\"\\\"}b2b,bCrxr?aab+b6bwobbOabb/byb5bYafbpu1bdbwbSazrkb8babmb5b=azv=awb6b*bNaEqgbJu1b?aPvgk\\\"\\\",2):f(\\\"\\\"}bdr*b/b0b\\\"\\\",2):f(\\\"\\\"}w7bfb\\\"\\\",2):f(\\\"\\\"{bXa=a@aybcbtbOa4bPa6pCaBvmbjbdbmbxbhbOaWaRawbbbBpSrCaQa1bPa0b\\\"\\\",2):f"));
$write("%s",("(\\\"\\\"{bjb.wZaYa,bwbZaXahw\\\"\\\",2):f(\\\"\\\"{b-bZa7b.bzrdb5pEakb+bew5bVagb=atb@rcbQqXa4b7b*bCa\\\"\\\",2):f(\\\"\\\"{j/bmbNazblb0bXa-b/bkbabcb7bBagbtk1bfbvbKvfvTaabdubu8sfb|o5klwwqtt-o1k2o\\\"\\\",2):f(\\\"\\\"}q\\\"\\\",2):f(\\\"\\\"{qQa|b/bUacbEa\\\"\\\",2):f(\\\"\\\"}bYaQa\\\"\\\",2):f(\\\"\\\"}bHjZtNaCagbtbxbWhmbwbXaDahr1bXaDpxbeb5bEatshtGaft<aubdb,bAtfbiv@pYa3b,byvfb/buvPaXabb1qxbgbkbmbPsjbWaCadbvb,b.blb,b,b0beb\\\"\\\",2):f(\\\"\\\"}bEatbgbubAaTa>a+bUubbhcCa,tOaab0btb7b9f*bXaBazb\\\"\\\",2):f(\\\"\\\"}b+bPaxbCaOawbzb<a2bYacb2bgb0bcb,b=aCaxb@aOa3bPa<skbFa?a/b-bRaUatbEa-b>smbgb\\\"\\\",2):f(\\\"\\\"}b8b0bHtPalbCr\\\"\\\",2):f(\\\"\\\"{bWa0btiOaAaFaZqabQa?a\\\"\\\",2):f(\\\"\\\"{bkbyb4bmbebgb,b6bTaUtWa|bCrbbzb8bFaibab4bCryblbTagbZbOrWa,bXq\\\"\\\",2):f(\\\"\\\"}bdb6byswbtsib+b,bdb8b.b2pXaEacb4b8bKidb/bSaCawb5bhbxbVa5b*dBaybDaVs|szs>r/k0o1o5k/o"));
$write("%s",("otzqot|q\\\"\\\",2):f(\\\"\\\"}o*qndQa7bus6issqs6ios@a/bPa*b\\\"\\\",2):f(\\\"\\\"}bwbBaQqOqwbHkVaUaTaBacbmb:pfbtb0b0bCr|bXaUaAaEjXambzb@a-bfb|b6b,b+b-bmbSrzbPqubTaVaBalr2bFaebybRaubzgeb6bdb5b7bHrnsCaCr-b3bUaCr7bRaXa,bSabbasAaNaYa/b@a.bcblb5b=r;r9rYqubjbcb9bzbjbRazb2bSceb7b2bQaZaCr@aGaqrmr\\\"\\\",2):f(\\\"\\\"{b/b5bOaubQa\\\"\\\",2):f(\\\"\\\"{b.bUaabwb1b/qkrir<aUavribTadbVajb,bIkWaBaFa-b\\\"\\\",2):f(\\\"\\\"{b7bPa,bWaxb6iqbRa1b-bab5bDaYaekDaUaPa7bDa@aFa1bSaEaFaMqKqvbAlmb7bNa1blbgbcbYaabPajb,q?ecbhbDaeqzb<qHpCpjb0pwb4plbYaZa-bibDaDa\\\"\\\",2):f(\\\"\\\"}b7b\\\"\\\",2):f(\\\"\\\"}bkbcbibjbRp5kxq+o3avq,o1kNm*o.o7btbbb|b2bIp;pBaDakb=ajbVjSaZaFaDa4bOp7bQaBaCpDafbBaFi\\\"\\\",2):f(\\\"\\\"{bcbwbebDaFaNaQa5bebUfkbdb+bib,bjbvb*b6bzb1babFa-pmbXaCaqpcbbbjbhbTaQa-bSa>aFa|b7bxbdbybHkeblbzb,bNa7bvbCaEahb<aCabb*bWhQaub*bWaQagbS"));
$write("%s",("a,bEa7b6bAaEamnMoxnmo8oJoPmao<nBo;amo=n?aEh6oloBo-bmnRnCa-arowbicmoZnko9oEaxnao5nXmBn0n.n/kLmMm1kKm|o9a|o|oul2kIm/b\\\"\\\",2):f(\\\"\\\"{f-aZhubeimoeopnjoWm9aEaQdSnZm3nXnXk:a-bao=aAa-aLnFnCaxnKn6l<a-b|eOnEnpn2n\\\"\\\",2):f(\\\"\\\"{nrnpnnn9nDn:aCa|e>n>aAa3nwnrn9aUmsnAaNlin|e1n4mmnznBa-aonhnfn*bvbtb/b-a+bIdantnbnkn@ainmnSe|egnln?aAaXm\\\"\\\",2):f(\\\"\\\"{bVmcnanFaYmWmUmHaSm9a|eTmxb8a+e-a1bUf8aPm1m8arb|e2b/k>m?m/k=m5k@m=kml:k7e8j6j|k1k;mBiBi3k/k8k*m6j6b-a+czbxbubHaqb6aqbSiTiRi5aqbebjj,bAfzb.bKfnb|fld6ixbEisfbgUkHhcjElsgCltcBa:jHl=kQlklBa?a:jvffi2g/h?aUhnlxkal?a>a:j6eZhrb3bglVhIhxlYgvl@aCa:j2b3bUiQfhk8fXk-bFk@a3aKa\\\"\\\",2):f(\\\"\\\"{b;a.b|bwbccIa3b1bpk,b|b0aYgel<k@hll>a@a:j.b?iVhsg?jZiblBarhggPcWk?ajiyk;k<jDa3a;d+cKfngbgfhubwb6i-aGkEk:a;bCk1b0b-b3a?a3akg6i.a:b:b,b?azk>jThwkBi6k4a4k"));
$write("%s",("/a0k;j4a-f.k-hCi9j5e7jmd*j0gVh|iaj=j;jZhwb+b-aPcdk/b8b1bPcxb;aQf-b:fZa\\\"\\\",2):f(\\\"\\\"{g|b.b5b-aVjKi3bIivb|bHjUi\\\"\\\",2):f(\\\"\\\"{gVf3bgf;a<b:b3b-a8b+bub,bxb2b2btb;aVhYgbj*i|i3arh5ani-jxb+j\\\"\\\",2):f(\\\"\\\"}jabVaTaRaOaHa6eEftiFfjb-agbebbbcbZaVa-abbVaEf-aZabbebSaHaebdb-aRhhbQabbZaVh@h7iPa8i,hnb-aSi/b3b4b.bHa8byb2b|b3btb2b-axb5b+b|hBi4awgyhVfTfMaFa=a|i-b*iIhiiGa+bJdwi9apg|fCcxbwb-bPaBaobThHfMa9aMaIa5axb3b.b4b0bxbzb-btbUfVhThjhMbub4b2bzb;azbLfccJa7b?a?aagIhCdYaOaVafbVaibNa=asg@h?a;a>a-aVaNaUawgYgvbpbEa|blgAaAa>aDa>anbJdubSczbJa2bIcag,fyfwfuf2bacYb-afgxc?aGaUe>a3a=gKaKa?angMbngGa>a:bngsbsg5ghgFgsbobsg*b-a4geg|fPgxbac1g\\\"\\\",2):f(\\\"\\\"}bnglg1aHg?abgrg\\\"\\\",2):f(\\\"\\\"{bHa2g0g-e:a:a\\\"\\\",2):f(\\\"\\\"}bHa@angJa\\\"\\\",2):f(\\\"\\\"}b5aAdteAangqgHa.bwbHa6a5bXf>azd:a,cNaXfwb.b;b/asg>ang-"));
$write("%s",("fag-a/b5a1aag2f7b-a@d-aQfybxcHa>a1aobob,c:a-a.b\\\"\\\",2):f(\\\"\\\"{bvbxb-a:b1d/b/a,fPcFf/b:b6aKa6e1b4eIa8\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"btb1b1bNaGatb5a+ctb,b-a\\\"\\\",2):f(\\\"\\\"{fyb3dMd-aDdBd@dmf/aob5a.d,d*d-b4b7eSc;axb+b.bbcZb0cbfJasdHa/aed+e0cGb/d,btb-b4aWbudpcgdLc=chchd6areOapc0cNb/a;bje/eGaHb5dedOb.a8aNd8aLdLa=a>aIaOaJapb6a+e5azb+cdcfbhc;aOaFdYd6aHaCa@aIaQd8aHa=a.cIbCbMd\\\"\\\",2):f(\\\"\\\"{cycvcocRapcXbocTa;b;bpbgbYdJaGbRanbQaJagbnbcb>dqc5dpbebnbOa8a0c4aJaTa5a+btb5bxbJaQa,c*cRa5a1bzc6aedMa0c3bldjd;aeded8ard5a6a5aedxb/btbvb2bxb,c1b4b3bxb1b0cocPa8aNapcMagdUc3b|b+b/b2b4arcFbnc4a=a?axbtc4aSbJcPbKckcic+bZb3b-bzcXbqcFb5aMa/ancvc+b+b|byb4a9cVbNa5aRb7cFbnbFbMapb2c.aMaFb.a4a5aJaOa-a-b|b-aeb5aicybHa<b/akc>a>aXb6aOb/a8a6a/apb4a1b.b3bvb4b1b3b2b-b.bvb4anb/aJaPa5a8a4a6apbEb5a5aBb,b9a4apbpbnb"));
$write("%s",("8anb4aGa=a:bJacb!\\\"\\\",2):f(\\\"\\\"})821(f\\\"\\\",2):f(\\\"\\\"{#~[2xha=s,y=z,23^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'Z3(yay,]99999[gnirtS wen=][c n3aea\\\"\\\",2):f(\\\"\\\"{)v]y3b&a(niam diov citats cilbup\\\"\\\",2):f(\\\"\\\"{RQ ssalc\\\"\\\",2):f(\\\"\\\"{4sfa cdlnl3c/a;maertStnirP/oi/avajL tuo/metsyS/gnal/avajn4bdateg@3doa2 kcats timil.v3dga]; V);R4aC3ecaL[c5aY4hha dohtem?3e;4nga repus&3ecaRQ@3cgassalc.=5koa(=:s;0=:c=:i;)\\\"\\\",2):f(\\\"\\\"}4ajaerudecorp03gqa(tnirp.biL.oken\\\"\\\",2):f(\\\"\\\"{/3bianoitcnufU6|sa(rtStup=niam^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9)"));
$write("%s",(":f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fla\\\"\\\",2):f(\\\"\\\"})36(f\\\"\\\",2):f(\\\"\\\"{#,43z3mba7D3a835oa(etirw.z;)tuo.N7aba(66b~auptuOPIZG.piz.litu.avaj wen=zv4,ka93623(f\\\"\\\",2):f(\\\"\\\"{#t:355aR0Z0Z/512152353/2/2166263=4/3141726??:1518191:1/n45da*6 L46ea1312~47\\\"\\\",2):f(\\\"\\\"{47fa41310?35Y9[83;M4dma(amirpmi oic$4[83jma++]371[]591[j55pani;RQ omtiroglaH35va;t:\\\"\\\",2):f(\\\"\\\"}%%%%\\\"\\\",2):f(\\\"\\\"}fi\\\"\\\",2):f(\\\"\\\"}*-84\\\"\\\",2):f(\\\"\\\"})867z3a(a]i[\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}+17\\\"\\\",2):f(\\\"\\\"{<84.;i:-i602\\\"\\\",2):f(\\\"\\\"{;i:911\\\"\\\",2):f(\\\"\\\"{;j:632|4,ea5526s@ajatnirP.tmfR@cfacnuf;P35datmf<36"));
$write("%s",("garopmi;PBagagakcapL3,ea3608#5dbapo5-?3cba-934jatnirp tesw:-ca69;;afantnirA5-ja9191(f\\\"\\\",2):f(\\\"\\\"{#f>31ca59$6awa,s(llAetirW;)(resUtxeT4Daca=:|5-ca38kAafanirp =33daS C;3-S=bca&(v43ba U4[U4qiaRQ margo#4/B3bjaS D : ; R*451B[83jL44qa. EPYT B C : ; A:5[83Cka)*,*(ETIRWD56haA B : ;A34ba [2c^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'47ia: ^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' ohce-A.ja(f\\\"\\\",2):f(\\\"\\"));
$write("%s",("\"{#(stupfEcdatniF3tca01z3sea%%%%:3[z3ipaparwyyon noitpoG3uw3Gca(n^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'Csba1p@a\\\"\\\",2):f(\\\"\\\"}7qba5nIa\\\"\\\",2):f(\\\"\\\"{aetirwf:oin\\\"\\\",2):f(\\\"\\\"})8(f\\\"\\\",2):f(\\\"\\\"{#>-)_(niamp3c*8nka(f\\\"\\\",2):f(\\\"\\\"{# cnirpOAoc8dma.OI[p]^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1"));
$write("%s",("^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'[06x#3cy4a\\\"\\\",2):f(\\\"\\\"}8cpadiov;oidts.dts vIaz5nV3d\\\"\\\",2):f(\\\"\\\"{3kkaenil-etirw64dva(,^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'s%^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'(gol.elosnoc;)^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f("));
$write("%s",("\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'73g\\\"\\\",2):f(\\\"\\\"}a^129^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' nioj.)1+n(yarrA>-)n(=fI3cwa^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"}54,1\\\"\\\",2):f(\\\"\\\"{.^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"# qes-er()|3cH3bba^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"p3lg3fw3hla1% ecalper.j4dea^128^I<c/arts(# pam(]Y"));
$write("%s",("ALPSID^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NOISIVID ERUDECORPA3cma.RQ .DI-MARGv3g53d|bNOITACIFITNEDI^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"[tac-yzal(s[qesod(^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))System.Console.Write($^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Put caffeine \\\"\\\",2):f(\\\"\\\"{(int)c\\\"\\\",2):f(\\\"\\\"} into the mixing bowl.^64^n^63^\\\"\\\",57):"));
$write("%s",("f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");M3pva^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Liquify contents ofE3oeaPour^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3w^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'4e\\\"\\\",2):f(\\\"\\\"{abaking dish.^64^n^64^nServes 164cma\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\"));
$write("%s",("\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}/****/e3a^15^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"),s[999999],*q=s;int main()\\\"\\\",2):f(\\\"\\\"{int n,m;for(;*p;)\\\"\\\",2):f(\\\"\\\"{n=(*p-5)%92+(p[1]-5)%92*87;p+=2;if(n>3999)for(m=(*p++-5)%92+6;m--;q++)*q=q[4000-n];else for(;n--;)*q++=*p++;\\\"\\\",2):f(\\\"\\\"}puts(s);return 0;\\\"\\\",2):f(\\\"\\\"}^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{s+=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(m=1;m<256;m*=2)s+=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f"));
$write("%s",("(\\\"\\\"\\\\\\\"\\\"00g,4,:^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+(c/m%2>0?^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4+^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\":^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")+^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\",^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";f(s);s=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4,:,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\"));
$write("%s",("\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";\\\"\\\",2):f(\\\"\\\"}f(s+s);for(c:Base64.getDecoder().decode(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"kaAREREX/I0ALn3n5ef6l/Pz8+fnz58/BOf5/7/hEX/OZzM5mCX/OczmZzBPn5+X/OczMznBL/nM5mZzBPu++fPPOc5zngnnOZzOZgnBMGAW7A==^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{c=c<0?256+c:c;for(i=0;i++<3;c/=8)f(c%8);f(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8*+8*+,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}f(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"@^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\"));
$write("%s",("\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");^1^\\\"\\\",4):f(\\\"\\\"'|sed -e^1^\\\"\\\",4):f(\\\"\\\"'s/^16^/^32^/g^1^\\\"\\\",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\\"'s/^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"/^16^q/g^1^\\\"\\\",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\\"'s/.*/print ^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^8^nquit/^1^\\\"\\\",4):f(\\\"\\\"'^3^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",2):f(\\\"\\\"}^1^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",4):f(\\\"\\\"');\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\""));
$write("%s",("\\\\\\\"\\\").split(\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",64):f(\\\"\\\"^\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");for(int i=1;i<a.length;a[0]+=a[i+1],i+=2)\\\"\\\",2):f(\\\"\\\"{a[0]+=\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",89):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".repeat(Integer.parseInt(a[i]));\\\"\\\",2):f(\\\"\\\"}System.out.print(a[0]);\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";FORiTO UPBtDO INTn:=ABSt[i];print(REPR(50+n%64)+c+REPR(50+n%8MOD8)+c+REPR(50+nMOD8)+b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"J\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+a)OD\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9)"));
$write("%s",(":f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"while(!=(S:length)0)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans c(S:read)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"D(c:to-integer)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 35 39\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 24 149\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"interp:library\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"afnix-sio\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans o(afnix:sio:OutputTerm)\\\"\\\",9):f(\\\"\\"));
$write("%s",("\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"o:write B\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");end;\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",1):f(\\\"\\\"nsys.exit 0'}\\\\\\\"\\\")\\\"\\\",0)]]></xsl:template></xsl:stylesheet>\\\":s.WriteByte(Asc(c)):Next:End Sub:End Module\")\nput=s\nprint\nqa!"));
end endmodule